library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

ENTITY FSM IS
	PORT(CLK,RST,RIGHT,LEFT, FLICK: IN STD_LOGIC;
		  LA,LB,LC,RA,RB,RC: OUT STD_LOGIC);
END ENTITY FSM;		  

ARCHITECTURE LOGIC OF FSM IS 

TYPE STATETYPE IS(I,L1,L2,L3,R1,R2,R3,F);
SIGNAL PRESENTS, NEXTS: STATETYPE;
BEGIN
	PROCESS(LEFT,RIGHT,PRESENTS)
	BEGIN
	CASE PRESENTS IS
	WHEN I=>
		IF(LEFT='1' AND RIGHT='1') THEN
			NEXTS<=F;
			ELSIF RIGHT='1' THEN
			NEXTS<=R1;
			ELSIF LEFT='1' THEN 
			NEXTS<=L1;
			ELSIF FLICK='1' THEN 
			NEXTS<=F;
			
			ELSE 
			NEXTS<=I;
			
			END IF;
			
	WHEN L1=>
			NEXTS<=L2;
	
	WHEN L2=>
			NEXTS<=L3;
	
	WHEN L3=>
			NEXTS<=I;

	WHEN R1=>
			NEXTS<=R2;
	
	WHEN R2=>
			NEXTS<=R3;		
	
	WHEN R3=>
			NEXTS<=I;
	WHEN F=>		
		IF(LEFT='1' AND RIGHT='1') THEN
			NEXTS<=F;
			ELSIF RIGHT='1' THEN
			NEXTS<=R1;
			ELSIF LEFT='1' THEN 
			NEXTS<=L1;
			ELSE NEXTS<=I;
			END IF;
	WHEN OTHERS=>
			nexts<=I;

	END CASE;
   END PROCESS;	
	
	PROCESS(CLK,RST)
	BEGIN
		IF RST='0' THEN
			PRESENTS<=I;
		ELSIF RISING_Edge(CLK) THEN
		PRESENTS<=NEXTS;
		END IF;
		END PROCESS;

		Lc<='1' WHEN (PRESENTS=L3 OR PRESENTS=F) ELSE '0';
		LB<='1' WHEN (PRESENTS=L3 OR PRESENTS=F OR PRESENTS=L2) ELSE '0';
		LA<='1' WHEN (PRESENTS=L3 OR PRESENTS=F OR PRESENTS=L1 OR PRESENTS=L2) ELSE '0';
		RA<='1' WHEN (PRESENTS=R3 OR PRESENTS=F OR PRESENTS=R1 OR PRESENTS=R2) ELSE '0';
		RB<='1' WHEN (PRESENTS=R2 OR PRESENTS=R3 OR PRESENTS=F) ELSE '0';
		RC<='1' WHEN (PRESENTS=R3 OR PRESENTS=F) ELSE '0';
END ARCHITECTURE LOGIC;

		